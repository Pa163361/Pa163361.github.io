magic
tech scmos
timestamp 1618808912
<< nwell >>
rect 0 0 24 20
<< ntransistor >>
rect 11 -16 13 -12
<< ptransistor >>
rect 11 6 13 14
<< ndiffusion >>
rect 10 -16 11 -12
rect 13 -16 14 -12
<< pdiffusion >>
rect 10 6 11 14
rect 13 6 14 14
<< ndcontact >>
rect 6 -16 10 -12
rect 14 -16 18 -12
<< pdcontact >>
rect 6 6 10 14
rect 14 6 18 14
<< polysilicon >>
rect 11 14 13 17
rect 11 -12 13 6
rect 11 -19 13 -16
<< polycontact >>
rect 7 -8 11 -4
<< metal1 >>
rect 0 22 24 26
rect 6 14 10 22
rect 14 -2 18 6
rect 2 -8 7 -4
rect 14 -6 24 -2
rect 14 -12 18 -6
rect 6 -20 10 -16
rect 6 -23 18 -20
<< labels >>
rlabel metal1 3 -7 4 -6 3 INP
rlabel metal1 17 -5 18 -4 1 Inv_out
rlabel metal1 14 -21 15 -20 1 gnd
rlabel metal1 11 23 12 24 5 vdd
<< end >>
