magic
tech scmos
timestamp 1619428530
<< ntransistor >>
rect 71 13 73 17
rect 79 13 81 17
<< ndiffusion >>
rect 70 13 71 17
rect 73 13 74 17
rect 78 13 79 17
rect 81 13 82 17
<< ndcontact >>
rect 66 13 70 17
rect 74 13 78 17
rect 82 13 86 17
<< polysilicon >>
rect 74 31 76 43
rect 71 29 76 31
rect 71 17 73 29
rect 79 17 81 52
rect 71 10 73 13
rect 79 10 81 13
<< polycontact >>
rect 75 47 79 51
rect 70 39 74 43
<< metal1 >>
rect 24 58 32 62
rect 56 58 91 62
rect 59 47 75 51
rect 59 28 63 47
rect 67 39 70 43
rect 67 36 72 39
rect 31 24 32 25
rect 56 24 63 28
rect 74 24 91 28
rect 58 16 66 21
rect 74 17 78 24
rect 62 13 66 16
rect 86 13 92 17
rect 87 12 92 13
rect 24 0 32 4
rect 56 0 91 4
<< m2contact >>
rect -1 23 4 28
rect 21 23 26 28
rect 31 25 36 30
rect 67 31 72 36
rect 53 16 58 21
rect 87 7 92 12
<< metal2 >>
rect 31 31 67 35
rect 31 30 36 31
rect -1 9 4 23
rect 21 21 26 23
rect 21 17 53 21
rect -1 7 87 9
rect -1 5 92 7
use inverter  inverter_0
timestamp 1618813994
transform 1 0 0 0 1 34
box 0 -34 24 28
use inverter  inverter_1
timestamp 1618813994
transform 1 0 32 0 1 34
box 0 -34 24 28
use inverter  inverter_2
timestamp 1618813994
transform 1 0 91 0 1 34
box 0 -34 24 28
use inverter  inverter_3
timestamp 1618813994
transform 1 0 115 0 1 34
box 0 -34 24 28
<< labels >>
rlabel metal1 86 24 88 28 7 XOR_out
rlabel polysilicon 72 27 73 28 1 B
rlabel polysilicon 80 40 81 41 1 B_bar
rlabel metal1 87 16 88 17 1 A
rlabel metal1 63 18 64 19 1 A_bar
<< end >>
