magic
tech scmos
timestamp 1618814130
use inverter  inverter_0
timestamp 1618813994
transform 1 0 0 0 1 34
box 0 -34 24 28
use inverter  inverter_1
timestamp 1618813994
transform 1 0 24 0 1 34
box 0 -34 24 28
<< end >>
