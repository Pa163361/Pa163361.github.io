* SPICE3 file created from or_five.ext - technology: scmos

.option scale=0.09u
.include TSMC_180nm.txt
.param SUPPLY=1.8
.global gnd vdd

Vol vdd gnd 'SUPPLY'

Vin_a A gnd pulse 0 1.8 0ps 1ps 1ps 10ns 20ns
Vin_b B gnd pulse 0 1.8 0ps 1ps 1ps 20ns 40ns
Vin_c C gnd pulse 0 1.8 0ps 1ps 1ps 40ns 80ns
Vin_d D gnd pulse 0 1.8 0ps 1ps 1ps 80ns 160ns
Vin_e E gnd pulse 0 1.8 0ps 1ps 1ps 160ns 320ns

M1000 or_five_output nor_five_output vdd vdd CMOSP w=8 l=2
+  ad=40 pd=26 as=80 ps=52
M1001 or_five_output nor_five_output gnd gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=88 ps=76
M1002 a_100_44# A vdd vdd CMOSP w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1003 a_108_44# B a_100_44# vdd CMOSP w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1004 a_116_44# C a_108_44# vdd CMOSP w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1005 a_124_44# D a_116_44# vdd CMOSP w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1006 nor_five_output E a_124_44# vdd CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1007 nor_five_output A gnd gnd CMOSN w=4 l=2
+  ad=68 pd=58 as=0 ps=0
M1008 gnd B nor_five_output gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 nor_five_output C gnd gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 gnd D nor_five_output gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 nor_five_output E gnd gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0

C0 nor_five_output or_five_output 0.1fF
C1 nor_five_output gnd 0.5fF
C2 vdd or_five_output 0.1fF
C3 or_five_output gnd 0.0fF
C4 vdd nor_five_output 0.1fF
C5 vdd vdd 0.1fF
C6 nor_five_output vdd 0.1fF
C7 vdd or_five_output 0.0fF
C8 gnd gnd 0.3fF
C9 or_five_output gnd 0.1fF
C10 vdd gnd 0.2fF
C11 nor_five_output gnd 0.9fF
C12 vdd gnd 2.0fF

.tran 0.1n 350n

.control

run

plot v(A) v(B) v(C) v(D) v(E)
plot v(or_five_output)

.endc

.end
