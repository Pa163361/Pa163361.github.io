* SPICE3 file created from or_three.ext - technology: scmos

.option scale=0.09u
.include TSMC_180nm.txt
.param SUPPLY=1.8
.global gnd vdd

Vdd vdd gnd 'SUPPLY'

Vin_a A gnd pulse 0 1.8 0ns 1ps 1ps 10ns 20ns
Vin_b B gnd pulse 0 1.8 0ns 1ps 1ps 20ns 40ns
Vin_c C gnd pulse 0 1.8 0ns 1ps 1ps 40ns 80ns

M1000 or_three_output NOR_three_out vdd vdd CMOSP w=8 l=2
+  ad=40 pd=26 as=80 ps=52
M1001 or_three_output NOR_three_out gnd gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=64 ps=56
M1002 a_108_44# A vdd vdd CMOSP w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1003 a_116_44# B a_108_44# vdd CMOSP w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1004 NOR_three_out C a_116_44# vdd CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1005 NOR_three_out A gnd gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=0 ps=0
M1006 gnd B NOR_three_out gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 NOR_three_out C gnd gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0

C0 vdd or_three_output 0.1fF
C1 NOR_three_out gnd 0.3fF
C2 vdd NOR_three_out 0.1fF
C3 or_three_output gnd 0.0fF
C4 vdd vdd 0.1fF
C5 NOR_three_out vdd 0.1fF
C6 vdd or_three_output 0.0fF
C7 NOR_three_out or_three_output 0.1fF
C8 gnd gnd 0.3fF
C9 or_three_output gnd 0.1fF
C10 vdd gnd 0.2fF
C11 NOR_three_out gnd 0.9fF
C12 vdd gnd 1.5fF

.tran 0.1n 200n

.control

run

plot v(A) v(B) v(C)
plot v(or_three_output)

.endc

.end
