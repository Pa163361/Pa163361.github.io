* SPICE3 file created from inverter.ext - technology: scmos

.option scale=0.09u
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.global gnd vdd

Vdd vdd gnd 'SUPPLY'

Vin INP gnd 0

M1000 Inv_out INP vdd vdd CMOSP w=8 l=2
+  ad=40 pd=26 as=40 ps=26
M1001 Inv_out INP gnd gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=20 ps=18

C0 INP Inv_out 0.1fF
C1 vdd Inv_out 0.1fF
C2 INP gnd 0.0fF
C3 Inv_out gnd 0.1fF
C4 INP vdd 0.1fF
C5 vdd vdd 0.0fF
C6 Inv_out vdd 0.0fF
C7 gnd gnd 0.1fF
C8 Inv_out gnd 0.1fF
C9 vdd gnd 0.1fF
C10 INP gnd 0.2fF
C11 vdd gnd 0.5fF

.tran 0.1n 200n

.control

run
plot v(Inv_out)

.endc

.end
