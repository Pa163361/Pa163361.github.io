* SPICE3 file created from xor_gate.ext - technology: scmos

.option scale=0.09u
.include TSMC_180nm.txt
.param SUPPLY=1.8
.global gnd vdd

Vdd vdd gnd 'SUPPLY'

Vin_a A gnd 1.8
Vin_a_bar A_bar gnd 0
Vin_b B gnd 0
Vin_b_bar B_bar gnd 1.8

M1000 final_out out_1 vdd vdd CMOSP w=8 l=2
+  ad=40 pd=26 as=160 ps=104
M1001 final_out out_1 gnd gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=80 ps=72
M1002 out_1 XOR_out vdd vdd CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1003 out_1 XOR_out gnd gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1004 B_bar B vdd vdd CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1005 B_bar B gnd gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1006 A_bar A vdd vdd CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1007 A_bar A gnd gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1008 XOR_out B A_bar gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=20 ps=18
M1009 A B_bar XOR_out gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
C0 out_1 XOR_out 0.1fF
C1 out_1 final_out 0.1fF
C2 A A 0.0fF
C3 gnd A 0.0fF
C4 vdd B 0.1fF
C5 vdd A 0.1fF
C6 vdd XOR_out 0.1fF
C7 vdd final_out 0.0fF
C8 B_bar B 0.1fF
C9 XOR_out A 0.1fF
C10 gnd XOR_out 0.0fF
C11 final_out gnd 0.0fF
C12 gnd A_bar 0.0fF
C13 vdd B_bar 0.0fF
C14 vdd A_bar 0.0fF
C15 vdd B_bar 0.2fF
C16 vdd vdd 0.0fF
C17 gnd B 0.0fF
C18 A A_bar 0.1fF
C19 vdd out_1 0.1fF
C20 gnd B_bar 0.0fF
C21 vdd vdd 0.1fF
C22 out_1 vdd 0.1fF
C23 vdd vdd 0.0fF
C24 B A_bar 0.1fF
C25 out_1 gnd 0.1fF
C26 XOR_out B_bar 0.1fF
C27 B_bar A_bar 0.0fF
C28 XOR_out A_bar 0.0fF
C29 vdd final_out 0.1fF
C30 A_bar A_bar 0.0fF
C31 vdd A_bar 0.1fF
C32 B B 0.0fF
C33 B B_bar 0.1fF
C34 A gnd 0.0fF
C35 A_bar gnd 0.0fF
C36 B gnd 0.2fF
C37 A_bar gnd 0.8fF
C38 A gnd 1.5fF
C39 vdd gnd 0.5fF
C40 B_bar gnd 0.5fF
C41 B gnd 0.7fF
C42 vdd gnd 0.5fF
C43 XOR_out gnd 0.3fF
C44 gnd gnd 0.6fF
C45 final_out gnd 0.1fF
C46 vdd gnd 0.5fF
C47 out_1 gnd 0.3fF
C48 vdd gnd 1.0fF

.tran 0.1n 200n

.control

run

plot v(A)
plot v(B)
plot v(final_out)

.endc

.end
