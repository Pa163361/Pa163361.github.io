magic
tech scmos
timestamp 1618810418
<< nwell >>
rect 0 0 32 20
<< ntransistor >>
rect 11 -26 13 -22
rect 19 -26 21 -22
<< ptransistor >>
rect 11 6 13 14
rect 19 6 21 14
<< ndiffusion >>
rect 10 -26 11 -22
rect 13 -26 19 -22
rect 21 -26 22 -22
<< pdiffusion >>
rect 10 6 11 14
rect 13 6 14 14
rect 18 6 19 14
rect 21 6 22 14
<< ndcontact >>
rect 6 -26 10 -22
rect 22 -26 26 -22
<< pdcontact >>
rect 6 6 10 14
rect 14 6 18 14
rect 22 6 26 14
<< polysilicon >>
rect 11 14 13 17
rect 19 14 21 17
rect 11 -22 13 6
rect 19 -1 21 6
rect 19 -3 24 -1
rect 22 -19 24 -3
rect 19 -21 24 -19
rect 19 -22 21 -21
rect 11 -29 13 -26
rect 19 -29 21 -26
<< polycontact >>
rect 7 -7 11 -3
rect 18 -15 22 -11
<< metal1 >>
rect -1 24 33 28
rect 6 14 10 24
rect 22 14 26 24
rect 14 -2 18 6
rect 3 -7 7 -3
rect 14 -6 30 -2
rect 26 -10 33 -6
rect 3 -15 18 -11
rect 26 -26 30 -10
rect 6 -30 10 -26
rect -1 -34 32 -30
<< labels >>
rlabel metal1 4 -5 5 -4 3 A
rlabel metal1 4 -12 5 -11 3 B
rlabel metal1 29 -9 30 -8 7 Out
rlabel pdcontact 6 6 10 14 1 pm_s_l
rlabel pdcontact 22 6 26 14 1 pm_s_r
rlabel metal1 17 -33 18 -32 1 Gnd
rlabel metal1 16 25 17 26 5 Vdd
<< end >>
