magic
tech scmos
timestamp 1619449071
<< nwell >>
rect 87 38 135 58
<< ntransistor >>
rect 98 8 100 12
rect 106 8 108 12
rect 114 8 116 12
rect 122 8 124 12
<< ptransistor >>
rect 98 44 100 52
rect 106 44 108 52
rect 114 44 116 52
rect 122 44 124 52
<< ndiffusion >>
rect 97 8 98 12
rect 100 8 101 12
rect 105 8 106 12
rect 108 8 109 12
rect 113 8 114 12
rect 116 8 117 12
rect 121 8 122 12
rect 124 8 125 12
<< pdiffusion >>
rect 97 44 98 52
rect 100 44 106 52
rect 108 44 114 52
rect 116 44 122 52
rect 124 44 125 52
<< ndcontact >>
rect 93 8 97 12
rect 101 8 105 12
rect 109 8 113 12
rect 117 8 121 12
rect 125 8 129 12
<< pdcontact >>
rect 93 44 97 52
rect 125 44 129 52
<< polysilicon >>
rect 98 52 100 55
rect 106 52 108 55
rect 114 52 116 55
rect 122 52 124 55
rect 98 43 100 44
rect 94 41 100 43
rect 94 15 96 41
rect 106 39 108 44
rect 104 37 108 39
rect 104 17 106 37
rect 104 15 108 17
rect 94 13 100 15
rect 98 12 100 13
rect 106 12 108 15
rect 114 12 116 44
rect 122 40 124 44
rect 122 38 126 40
rect 124 17 126 38
rect 122 15 126 17
rect 122 12 124 15
rect 98 5 100 8
rect 106 5 108 8
rect 114 5 116 8
rect 122 5 124 8
<< polycontact >>
rect 90 33 94 37
rect 100 33 104 37
rect 110 29 114 33
rect 120 29 124 33
<< metal1 >>
rect 87 58 135 62
rect 93 52 97 58
rect 129 28 133 52
rect 129 24 136 28
rect 129 19 133 24
rect 101 15 133 19
rect 101 12 105 15
rect 117 12 121 15
rect 93 4 97 8
rect 109 4 113 8
rect 125 4 129 8
rect 87 0 135 4
use inverter  inverter_0
timestamp 1618813994
transform 1 0 135 0 1 34
box 0 -34 24 28
<< labels >>
rlabel metal1 110 59 111 60 5 vdd
rlabel metal1 109 1 110 2 1 gnd
rlabel polysilicon 95 35 96 36 1 A
rlabel polysilicon 105 36 106 37 1 B
rlabel polysilicon 114 36 115 37 1 C
rlabel polysilicon 124 26 125 27 1 D
<< end >>
