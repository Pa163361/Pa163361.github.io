* SPICE3 file created from and_gate.ext - technology: scmos

.option scale=0.09u
.include TSMC_180nm.txt
.param SUPPLY=1.8
.global gnd vdd

Vdd vdd gnd 'SUPPLY'

Vin_a A gnd 1.8
Vin_b B gnd 0

M1000 Inv_out Out vdd vdd CMOSP w=8 l=2
+  ad=40 pd=26 as=120 ps=78
M1001 Inv_out Out gnd gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1002 Out A vdd vdd CMOSP w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1003 vdd B Out vdd CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 C A gnd gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1005 Out B C gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
C0 Inv_out gnd 0.0fF
C1 Out gnd 0.1fF
C2 vdd Inv_out 0.0fF
C3 Out Inv_out 0.1fF
C4 vdd Out 0.1fF
C5 vdd Inv_out 0.1fF
C6 vdd vdd 0.1fF
C7 Out vdd 0.2fF
C8 gnd gnd 0.3fF
C9 Inv_out gnd 0.1fF
C10 vdd gnd 0.2fF
C11 Out gnd 0.6fF
C12 vdd gnd 1.3fF

.tran 0.1n 200n

.control

run

plot v(Inv_out)

.endc

.end
