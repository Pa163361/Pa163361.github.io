magic
tech scmos
timestamp 1619431676
<< nwell >>
rect 80 38 128 58
<< ntransistor >>
rect 91 8 93 12
rect 99 8 101 12
rect 107 8 109 12
rect 115 8 117 12
<< ptransistor >>
rect 91 44 93 52
rect 99 44 101 52
rect 107 44 109 52
rect 115 44 117 52
<< ndiffusion >>
rect 90 8 91 12
rect 93 8 99 12
rect 101 8 107 12
rect 109 8 115 12
rect 117 8 118 12
<< pdiffusion >>
rect 90 44 91 52
rect 93 44 94 52
rect 98 44 99 52
rect 101 44 102 52
rect 106 44 107 52
rect 109 44 110 52
rect 114 44 115 52
rect 117 44 118 52
<< ndcontact >>
rect 86 8 90 12
rect 118 8 122 12
<< pdcontact >>
rect 86 44 90 52
rect 94 44 98 52
rect 102 44 106 52
rect 110 44 114 52
rect 118 44 122 52
<< polysilicon >>
rect 91 52 93 55
rect 99 52 101 55
rect 107 52 109 55
rect 115 52 117 55
rect 91 43 93 44
rect 87 41 93 43
rect 87 16 89 41
rect 99 37 101 44
rect 98 35 101 37
rect 107 38 109 44
rect 115 38 117 44
rect 107 36 111 38
rect 115 36 121 38
rect 98 24 100 35
rect 96 22 100 24
rect 87 14 93 16
rect 91 12 93 14
rect 96 15 98 22
rect 109 16 111 36
rect 119 16 121 36
rect 96 13 101 15
rect 99 12 101 13
rect 107 14 111 16
rect 115 14 121 16
rect 107 12 109 14
rect 115 12 117 14
rect 91 5 93 8
rect 99 5 101 8
rect 107 5 109 8
rect 115 5 117 8
<< polycontact >>
rect 83 33 87 37
rect 94 30 98 34
rect 105 28 109 32
rect 115 28 119 32
<< metal1 >>
rect 80 58 128 62
rect 86 52 90 58
rect 102 52 106 58
rect 118 52 122 58
rect 94 41 98 44
rect 110 41 114 44
rect 94 37 126 41
rect 122 28 126 37
rect 122 24 128 28
rect 122 8 126 24
rect 86 4 90 8
rect 80 0 128 4
use inverter  inverter_0
timestamp 1618813994
transform 1 0 128 0 1 34
box 0 -34 24 28
<< labels >>
rlabel metal1 103 59 104 60 5 vdd
rlabel metal1 99 1 100 2 1 gnd
rlabel metal1 125 26 126 27 7 nand_three_out
rlabel polysilicon 87 33 88 34 1 A
rlabel polysilicon 98 31 99 32 1 B
rlabel polysilicon 109 30 110 31 1 C
rlabel polysilicon 119 31 120 32 1 D
<< end >>
