magic
tech scmos
timestamp 1618813994
<< nwell >>
rect 0 0 24 20
<< ntransistor >>
rect 11 -20 13 -16
<< ptransistor >>
rect 11 6 13 14
<< ndiffusion >>
rect 10 -20 11 -16
rect 13 -20 14 -16
<< pdiffusion >>
rect 10 6 11 14
rect 13 6 14 14
<< ndcontact >>
rect 6 -20 10 -16
rect 14 -20 18 -16
<< pdcontact >>
rect 6 6 10 14
rect 14 6 18 14
<< polysilicon >>
rect 11 14 13 17
rect 11 -16 13 6
rect 11 -23 13 -20
<< polycontact >>
rect 7 -10 11 -6
<< metal1 >>
rect 0 24 24 28
rect 6 14 10 24
rect 14 -6 18 6
rect 0 -10 7 -6
rect 14 -10 24 -6
rect 14 -16 18 -10
rect 6 -30 10 -20
rect 0 -34 24 -30
<< labels >>
rlabel metal1 3 -9 4 -8 3 INP
rlabel metal1 14 -31 15 -30 1 gnd
rlabel metal1 13 25 14 26 5 vdd
rlabel metal1 17 -9 18 -8 1 Inv_out
<< end >>
