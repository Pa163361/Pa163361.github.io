magic
tech scmos
timestamp 1618810167
use nand_two  nand_two_0
timestamp 1618801919
transform 1 0 0 0 1 34
box 0 -34 32 28
<< end >>
