* SPICE3 file created from or_gate.ext - technology: scmos

.option scale=0.09u
.include TSMC_180nm.txt
.param SUPPLY=1.8
.global gnd vdd

Vdd vdd gnd 'SUPPLY'

Vin_a A gnd 1.8
Vin_a_bar A_bar gnd 0
Vin_b B gnd 0
Vin_b_bar B_bar gnd 1.8

M1000 or_gate_output or_out vdd vdd CMOSP w=8 l=2
+  ad=40 pd=26 as=80 ps=52
M1001 or_gate_output or_out gnd gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=60 ps=54
M1002 C B vdd vdd CMOSP w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1003 or_out A C vdd CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1004 or_out B gnd gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1005 gnd A or_out gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
C0 or_out gnd 0.2fF
C1 vdd vdd 0.1fF
C2 vdd or_out 0.1fF
C3 or_gate_output gnd 0.0fF
C4 vdd or_gate_output 0.1fF
C5 vdd or_gate_output 0.0fF
C6 or_out or_gate_output 0.1fF
C7 gnd gnd 0.3fF
C8 or_gate_output gnd 0.1fF
C9 vdd gnd 0.2fF
C10 or_out gnd 0.4fF
C11 vdd gnd 1.3fF

.tran 01.n 200n

.control

run

plot v(A)
plot v(B)
plot v(or_gate_output)

.endc

.end
