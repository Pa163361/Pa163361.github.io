* SPICE3 file created from and_four.ext - technology: scmos

.option scale=0.09u
.include TSMC_180nm.txt
.param SUPPLY=1.8
.global gnd vdd

Vdd vdd gnd 'SUPPLY'

Vin_a A gnd pulse 0 1.8 0ns 1ps 1ps 10ns 20ns
Vin_b B gnd pulse 0 1.8 0ns 1ps 1ps 20ns 40ns
Vin_c C gnd pulse 0 1.8 0ns 1ps 1ps 40ns 80ns
Vin_d D gnd pulse 0 1.8 0ns 1ps 1ps 80ns 160ns

M1000 and_four_output nand_three_out vdd vdd CMOSP w=8 l=2
+  ad=40 pd=26 as=168 ps=106
M1001 and_four_output nand_three_out gnd gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1002 nand_three_out A vdd vdd CMOSP w=8 l=2
+  ad=96 pd=56 as=0 ps=0
M1003 vdd B nand_three_out vdd CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 nand_three_out C vdd vdd CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 vdd D nand_three_out vdd CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 a_93_8# A gnd gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1007 a_101_8# B a_93_8# gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1008 a_109_8# C a_101_8# gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1009 nand_three_out D a_109_8# gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0

C0 vdd vdd 0.2fF
C1 nand_three_out vdd 0.5fF
C2 vdd and_four_output 0.0fF
C3 nand_three_out and_four_output 0.1fF
C4 nand_three_out gnd 0.1fF
C5 vdd and_four_output 0.1fF
C6 and_four_output gnd 0.0fF
C7 vdd nand_three_out 0.1fF
C8 a_109_8# gnd 0.0fF
C9 a_101_8# gnd 0.0fF
C10 a_93_8# gnd 0.0fF
C11 gnd gnd 0.4fF
C12 and_four_output gnd 0.1fF
C13 vdd gnd 0.2fF
C14 nand_three_out gnd 0.9fF
C15 vdd gnd 1.7fF

.tran 0.1n 200n

.control

run

plot v(A)
plot v(B)
plot v(C)
plot v(D)
plot v(and_four_output)

.endc

.end
